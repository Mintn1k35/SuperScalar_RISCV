
module LSU(
	// Input signals
		


	// Output signals	
);
endmodule: LSU






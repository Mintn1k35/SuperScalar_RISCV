`timescale 1ns/1ps

`include "../rtl/name.v"

module tb_name;

	// Input signals
	

	// Output signals
	


	initial begin
		$dumpfile("wave_file/tb_name.vcd");
		$dumpvars(0, tb_name);
	end

	
	initial begin

	end


	name name_instance();
endmodule

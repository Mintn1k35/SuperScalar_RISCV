
`include "define_module.v"
module AU(
	// Input signals
	


	// Output signals	
);
endmodule






`include "Cache_Controller"
module Core(
	// Input signals
	


	// Output signals	
);
endmodule: Core






module name(
	// Input signals
	


	// Output signals	
);
endmodule





